library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package network_types is
    type mem is array (natural range <>) of std_logic_vector;
    
end package network_types;